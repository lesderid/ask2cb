/*
两个2位二进制数的乘法，结果输出到数码管显示
*/
module mlt(a,b,c,en);

input[1:0] a,b;
output[7:0] c;
reg[7:0] c;
output en;

wire[3:0] c_tmp;

assign en=0;
assign c_tmp=a*b;

always@(c_tmp)
begin
	case(c_tmp)
		4'b0000:
			c=8'b0000_0011;
		4'b0001:
			c=8'b1001_1111;
		4'b0010:
			c=8'b0010_0101;
		4'b0011:
			c=8'b0000_1101;
		4'b0100:
			c=8'b1001_1001;
		4'b0101:
			c=8'b0100_1001;
		4'b0110:
			c=8'b0100_0001;
		4'b0111:
			c=8'b0001_1111;
		4'b1000:
			c=8'b0000_0001;
		4'b1001:
			c=8'b0001_1001;
		4'b1010:
			c=8'b0001_0001;
		4'b1011:
			c=8'b1100_0001;
		4'b1100:
			c=8'b0110_0011;
		4'b1101:
			c=8'b1000_0101;
		4'b1110:
			c=8'b0110_0001;
		4'b1111:
			c=8'b0111_0001;
	 endcase
end
endmodule 