LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.ALL;
USE  IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY  beep1 IS
  PORT(
        CLK:IN STD_LOGIC;
      --  DIGIT:BUFFER STD_LOGIC_VECTOR(6 DOWNTO 0);
        SPEAKER	:OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE SONG OF beep1 IS
SIGNAL DRIVER,ORIGIN:STD_LOGIC_VECTOR(12 DOWNTO 0);
SIGNAL COUNTER:INTEGER RANGE 0 TO 140;
SIGNAL COUNTER1:INTEGER RANGE 0 TO 3;
SIGNAL COUNTER2:INTEGER RANGE 1 TO 10000000;
SIGNAL DIGIT  :STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL COUNT  :STD_LOGIC_VECTOR(1 DOWNTO 0); 
SIGNAL CARRIER,CLK_4MHZ,CLK_4HZ:STD_LOGIC;
  BEGIN
PROCESS(CLK)
BEGIN
IF CLK'EVENT AND CLK='1' THEN
   IF COUNTER1=1 THEN CLK_4MHZ<='1';
      COUNTER1<=2;
   ELSIF COUNTER1=3 THEN CLK_4MHZ<='0';
      COUNTER1<=0;
   ELSE COUNTER1<=COUNTER1+1;
   END IF;
   
   IF COUNTER2=5000000 THEN CLK_4HZ<='1';
      COUNTER2<=5000001;
   ELSIF COUNTER2=10000000 THEN CLK_4HZ<='0';
      COUNTER2<=1;
   ELSE COUNTER2<=COUNTER2+1;
   END IF;
END IF;
END PROCESS;

PROCESS(CLK_4MHZ)
BEGIN
 IF CLK_4MHZ'EVENT AND CLK_4MHZ='1' THEN
    IF DRIVER="1111111111111"THEN
       CARRIER<='1';
       DRIVER<=ORIGIN;
ELSE
DRIVER<=DRIVER+1;
CARRIER<='0';
END IF;
END IF;
END PROCESS;

PROCESS(CARRIER)
BEGIN
IF CARRIER'EVENT AND CARRIER='1' THEN
COUNT<=COUNT+1;
IF COUNT="00"THEN
SPEAKER<='1';
ELSE
SPEAKER<='0';
END IF;
END IF;
END PROCESS;

PROCESS(CLK_4HZ)
BEGIN
IF CLK_4HZ'EVENT AND CLK_4HZ='1' THEN
 IF COUNTER=140 THEN
COUNTER<=0;
ELSE COUNTER<=COUNTER+1;
END IF;
END IF;
CASE COUNTER IS
WHEN 0  =>DIGIT<="0000011";          WHEN 1  =>DIGIT<="0000011";
WHEN 2  =>DIGIT<="0000011";          WHEN 3  =>DIGIT<="0000011";
WHEN 4  =>DIGIT<="0000101";          WHEN 5  =>DIGIT<="0000101";
WHEN 6  =>DIGIT<="0000101";          WHEN 7  =>DIGIT<="0000110";
WHEN 8  =>DIGIT<="0001000";          WHEN 9  =>DIGIT<="0001000";
WHEN 10 =>DIGIT<="0001000";          WHEN 11 =>DIGIT<="0010000";
WHEN 12 =>DIGIT<="0000110";          WHEN 13 =>DIGIT<="0001000";
WHEN 14 =>DIGIT<="0000101";          WHEN 15 =>DIGIT<="0000101";
WHEN 16 =>DIGIT<="0101000";          WHEN 17 =>DIGIT<="0101000";
WHEN 18 =>DIGIT<="0101000";          WHEN 19 =>DIGIT<="1000000";
WHEN 20 =>DIGIT<="0110000";          WHEN 21 =>DIGIT<="0101000";
WHEN 22 =>DIGIT<="0011000";          WHEN 23 =>DIGIT<="0101000";
WHEN 24 =>DIGIT<="0010000";          WHEN 25 =>DIGIT<="0010000";
WHEN 26 =>DIGIT<="0010000";          WHEN 27 =>DIGIT<="0010000";
WHEN 28 =>DIGIT<="0010000";          WHEN 29 =>DIGIT<="0010000";
WHEN 30 =>DIGIT<="0000011";          WHEN 31 =>DIGIT<="0000000";
WHEN 32 =>DIGIT<="0010000";          WHEN 33 =>DIGIT<="0010000";
WHEN 34 =>DIGIT<="0010000";          WHEN 35 =>DIGIT<="0011000";
WHEN 36 =>DIGIT<="0000111";          WHEN 37 =>DIGIT<="0000111";
WHEN 38 =>DIGIT<="0000110";          WHEN 39 =>DIGIT<="0000110";
WHEN 40 =>DIGIT<="0000101";          WHEN 41 =>DIGIT<="0000101";
WHEN 42 =>DIGIT<="0000101";          WHEN 43 =>DIGIT<="0000110";
WHEN 44 =>DIGIT<="0001000";          WHEN 45 =>DIGIT<="0001000";
WHEN 46 =>DIGIT<="0010000";          WHEN 47 =>DIGIT<="0010000";
WHEN 48 =>DIGIT<="0000011";          WHEN 49 =>DIGIT<="0000011";
WHEN 50 =>DIGIT<="0001000";          WHEN 51 =>DIGIT<="0001000";
WHEN 52 =>DIGIT<="0000110";          WHEN 53 =>DIGIT<="0000101";
WHEN 54 =>DIGIT<="0000110";          WHEN 55 =>DIGIT<="0001000";
WHEN 56 =>DIGIT<="0000101";          WHEN 57 =>DIGIT<="0000101";
WHEN 58 =>DIGIT<="0000101";          WHEN 59 =>DIGIT<="0000101";
WHEN 60 =>DIGIT<="0000101";          WHEN 61 =>DIGIT<="0000101";
WHEN 62 =>DIGIT<="0000101";          WHEN 63 =>DIGIT<="0000101";
WHEN 64 =>DIGIT<="0011000";          WHEN 65 =>DIGIT<="0011000";
WHEN 66 =>DIGIT<="0011000";          WHEN 67 =>DIGIT<="0101000";
WHEN 68 =>DIGIT<="0000111";          WHEN 69 =>DIGIT<="0000111";
WHEN 70 =>DIGIT<="0010000";          WHEN 71 =>DIGIT<="0010000";
WHEN 72 =>DIGIT<="0000110";          WHEN 73 =>DIGIT<="0001000";
WHEN 74 =>DIGIT<="0000101";          WHEN 75 =>DIGIT<="0000101";
WHEN 76 =>DIGIT<="0000101";          WHEN 77 =>DIGIT<="0000101";
WHEN 78 =>DIGIT<="0000101";          WHEN 79 =>DIGIT<="0000101";
WHEN 80 =>DIGIT<="0000011";          WHEN 81 =>DIGIT<="0000101";
WHEN 82 =>DIGIT<="0000011";          WHEN 83 =>DIGIT<="0000011";
WHEN 84 =>DIGIT<="0000101";          WHEN 85 =>DIGIT<="0000110";
WHEN 86 =>DIGIT<="0000111";          WHEN 87 =>DIGIT<="0010000";
WHEN 88 =>DIGIT<="0000110";          WHEN 89 =>DIGIT<="0000110";
WHEN 90 =>DIGIT<="0000110";          WHEN 91 =>DIGIT<="0000110";
WHEN 92 =>DIGIT<="0000110";          WHEN 93 =>DIGIT<="0000110";
WHEN 94 =>DIGIT<="0000101";          WHEN 95 =>DIGIT<="0000110";
WHEN 96 =>DIGIT<="0001000";          WHEN 97 =>DIGIT<="0001000";
WHEN 98 =>DIGIT<="0001000";          WHEN 99 =>DIGIT<="0010000";
WHEN 100=>DIGIT<="0101000";          WHEN 101=>DIGIT<="0101000";
WHEN 102=>DIGIT<="0101000";          WHEN 103=>DIGIT<="0011000";
WHEN 104=>DIGIT<="0010000";          WHEN 105=>DIGIT<="0010000";
WHEN 106=>DIGIT<="0011000";          WHEN 107=>DIGIT<="0010000";
WHEN 108=>DIGIT<="0001000";          WHEN 109=>DIGIT<="0001000";
WHEN 110=>DIGIT<="0000110";          WHEN 111=>DIGIT<="0000101";
WHEN 112=>DIGIT<="0000011";          WHEN 113=>DIGIT<="0000011";
WHEN 114=>DIGIT<="0000011";          WHEN 115=>DIGIT<="0000011";
WHEN 116=>DIGIT<="0001000";          WHEN 117=>DIGIT<="0001000";
WHEN 118=>DIGIT<="0000110";          WHEN 119=>DIGIT<="0001000";
WHEN 120=>DIGIT<="0000110";          WHEN 121=>DIGIT<="0000011";
WHEN 122=>DIGIT<="0000011";          WHEN 123=>DIGIT<="0010000";
WHEN 124=>DIGIT<="0000011";          WHEN 125=>DIGIT<="0000101";
WHEN 126=>DIGIT<="0000110";          WHEN 127=>DIGIT<="0001000";
WHEN 128=>DIGIT<="0000101";          WHEN 129=>DIGIT<="0000101";
WHEN 130=>DIGIT<="0000101";          WHEN 131=>DIGIT<="0000101";
WHEN 132=>DIGIT<="0000101";          WHEN 133=>DIGIT<="0000101";
WHEN 134=>DIGIT<="0000101";          WHEN 135=>DIGIT<="0000101";
WHEN 136=>DIGIT<="0000000";          WHEN 137=>DIGIT<="0000000";
WHEN 138=>DIGIT<="0000000";          WHEN 139=>DIGIT<="0000000";
WHEN OTHERS=>DIGIT<="0000000";
END CASE;
CASE DIGIT IS
  WHEN "0000011"=>ORIGIN<="0100001001100";
  WHEN "0000101"=>ORIGIN<="0110000010001";
  WHEN "0000110"=>ORIGIN<="0111000111110";
  WHEN "0000111"=>ORIGIN<="1000000101101";
  WHEN "0001000"=>ORIGIN<="1000100010001";
  WHEN "0010000"=>ORIGIN<="1001010110010";
  WHEN "0011000"=>ORIGIN<="1010000100101";
  WHEN "0101000"=>ORIGIN<="1011000001000";
  WHEN "0110000"=>ORIGIN<="1011100011110";
  WHEN "1000000"=>ORIGIN<="1100010001000";
WHEN OTHERS=>ORIGIN<="1111111111111";
END CASE;
END PROCESS;
END SONG;




